----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 14.10.2018 09:15:59
-- Design Name: 
-- Module Name: sigmoid_lut - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sigmoid_lut is
    Port ( clk : in STD_LOGIC;
           en : in STD_LOGIC;
           din : in STD_LOGIC_VECTOR (15 downto 0);
           dout : out STD_LOGIC_VECTOR (15 downto 0));
end sigmoid_lut;

architecture Behavioral of sigmoid_lut is
    type SIGMOID_LUT_TYPE is ARRAY(8191 downto 0) of STD_LOGIC_VECTOR(15 downto 0);
    signal lut : SIGMOID_LUT_TYPE := (x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FF", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FE", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FD", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FC", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FB", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00FA", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F9", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F8", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F7", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F6", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F5", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F4", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F3", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F2", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F1", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00F0", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EF", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00EE", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00ED", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EC", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EB", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00EA", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E9", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E8", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E7", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E6", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E5", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E4", x"00E3", x"00E3", x"00E3", x"00E3", x"00E3", x"00E3", x"00E3", x"00E3", x"00E3", x"00E3", x"00E2", x"00E2", x"00E2", x"00E2", x"00E2", x"00E2", x"00E2", x"00E2", x"00E2", x"00E2", x"00E1", x"00E1", x"00E1", x"00E1", x"00E1", x"00E1", x"00E1", x"00E1", x"00E1", x"00E0", x"00E0", x"00E0", x"00E0", x"00E0", x"00E0", x"00E0", x"00E0", x"00E0", x"00DF", x"00DF", x"00DF", x"00DF", x"00DF", x"00DF", x"00DF", x"00DF", x"00DF", x"00DE", x"00DE", x"00DE", x"00DE", x"00DE", x"00DE", x"00DE", x"00DE", x"00DE", x"00DD", x"00DD", x"00DD", x"00DD", x"00DD", x"00DD", x"00DD", x"00DD", x"00DD", x"00DC", x"00DC", x"00DC", x"00DC", x"00DC", x"00DC", x"00DC", x"00DC", x"00DB", x"00DB", x"00DB", x"00DB", x"00DB", x"00DB", x"00DB", x"00DB", x"00DA", x"00DA", x"00DA", x"00DA", x"00DA", x"00DA", x"00DA", x"00DA", x"00D9", x"00D9", x"00D9", x"00D9", x"00D9", x"00D9", x"00D9", x"00D9", x"00D8", x"00D8", x"00D8", x"00D8", x"00D8", x"00D8", x"00D8", x"00D8", x"00D7", x"00D7", x"00D7", x"00D7", x"00D7", x"00D7", x"00D7", x"00D6", x"00D6", x"00D6", x"00D6", x"00D6", x"00D6", x"00D6", x"00D6", x"00D5", x"00D5", x"00D5", x"00D5", x"00D5", x"00D5", x"00D5", x"00D4", x"00D4", x"00D4", x"00D4", x"00D4", x"00D4", x"00D4", x"00D3", x"00D3", x"00D3", x"00D3", x"00D3", x"00D3", x"00D3", x"00D2", x"00D2", x"00D2", x"00D2", x"00D2", x"00D2", x"00D2", x"00D1", x"00D1", x"00D1", x"00D1", x"00D1", x"00D1", x"00D1", x"00D0", x"00D0", x"00D0", x"00D0", x"00D0", x"00D0", x"00CF", x"00CF", x"00CF", x"00CF", x"00CF", x"00CF", x"00CF", x"00CE", x"00CE", x"00CE", x"00CE", x"00CE", x"00CE", x"00CD", x"00CD", x"00CD", x"00CD", x"00CD", x"00CD", x"00CC", x"00CC", x"00CC", x"00CC", x"00CC", x"00CC", x"00CC", x"00CB", x"00CB", x"00CB", x"00CB", x"00CB", x"00CB", x"00CA", x"00CA", x"00CA", x"00CA", x"00CA", x"00CA", x"00C9", x"00C9", x"00C9", x"00C9", x"00C9", x"00C9", x"00C8", x"00C8", x"00C8", x"00C8", x"00C8", x"00C8", x"00C7", x"00C7", x"00C7", x"00C7", x"00C7", x"00C6", x"00C6", x"00C6", x"00C6", x"00C6", x"00C6", x"00C5", x"00C5", x"00C5", x"00C5", x"00C5", x"00C5", x"00C4", x"00C4", x"00C4", x"00C4", x"00C4", x"00C3", x"00C3", x"00C3", x"00C3", x"00C3", x"00C3", x"00C2", x"00C2", x"00C2", x"00C2", x"00C2", x"00C1", x"00C1", x"00C1", x"00C1", x"00C1", x"00C1", x"00C0", x"00C0", x"00C0", x"00C0", x"00C0", x"00BF", x"00BF", x"00BF", x"00BF", x"00BF", x"00BF", x"00BE", x"00BE", x"00BE", x"00BE", x"00BE", x"00BD", x"00BD", x"00BD", x"00BD", x"00BD", x"00BC", x"00BC", x"00BC", x"00BC", x"00BC", x"00BB", x"00BB", x"00BB", x"00BB", x"00BB", x"00BA", x"00BA", x"00BA", x"00BA", x"00BA", x"00B9", x"00B9", x"00B9", x"00B9", x"00B9", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8", x"00B7", x"00B7", x"00B7", x"00B7", x"00B7", x"00B6", x"00B6", x"00B6", x"00B6", x"00B6", x"00B5", x"00B5", x"00B5", x"00B5", x"00B5", x"00B4", x"00B4", x"00B4", x"00B4", x"00B4", x"00B3", x"00B3", x"00B3", x"00B3", x"00B3", x"00B2", x"00B2", x"00B2", x"00B2", x"00B1", x"00B1", x"00B1", x"00B1", x"00B1", x"00B0", x"00B0", x"00B0", x"00B0", x"00B0", x"00AF", x"00AF", x"00AF", x"00AF", x"00AE", x"00AE", x"00AE", x"00AE", x"00AE", x"00AD", x"00AD", x"00AD", x"00AD", x"00AC", x"00AC", x"00AC", x"00AC", x"00AC", x"00AB", x"00AB", x"00AB", x"00AB", x"00AB", x"00AA", x"00AA", x"00AA", x"00AA", x"00A9", x"00A9", x"00A9", x"00A9", x"00A9", x"00A8", x"00A8", x"00A8", x"00A8", x"00A7", x"00A7", x"00A7", x"00A7", x"00A6", x"00A6", x"00A6", x"00A6", x"00A6", x"00A5", x"00A5", x"00A5", x"00A5", x"00A4", x"00A4", x"00A4", x"00A4", x"00A4", x"00A3", x"00A3", x"00A3", x"00A3", x"00A2", x"00A2", x"00A2", x"00A2", x"00A1", x"00A1", x"00A1", x"00A1", x"00A0", x"00A0", x"00A0", x"00A0", x"00A0", x"009F", x"009F", x"009F", x"009F", x"009E", x"009E", x"009E", x"009E", x"009D", x"009D", x"009D", x"009D", x"009C", x"009C", x"009C", x"009C", x"009C", x"009B", x"009B", x"009B", x"009B", x"009A", x"009A", x"009A", x"009A", x"0099", x"0099", x"0099", x"0099", x"0098", x"0098", x"0098", x"0098", x"0097", x"0097", x"0097", x"0097", x"0096", x"0096", x"0096", x"0096", x"0096", x"0095", x"0095", x"0095", x"0095", x"0094", x"0094", x"0094", x"0094", x"0093", x"0093", x"0093", x"0093", x"0092", x"0092", x"0092", x"0092", x"0091", x"0091", x"0091", x"0091", x"0090", x"0090", x"0090", x"0090", x"008F", x"008F", x"008F", x"008F", x"008E", x"008E", x"008E", x"008E", x"008D", x"008D", x"008D", x"008D", x"008C", x"008C", x"008C", x"008C", x"008B", x"008B", x"008B", x"008B", x"008A", x"008A", x"008A", x"008A", x"0089", x"0089", x"0089", x"0089", x"0088", x"0088", x"0088", x"0088", x"0087", x"0087", x"0087", x"0087", x"0086", x"0086", x"0086", x"0086", x"0085", x"0085", x"0085", x"0085", x"0084", x"0084", x"0084", x"0084", x"0083", x"0083", x"0083", x"0083", x"0082", x"0082", x"0082", x"0082", x"0081", x"0081", x"0081", x"0081", x"0080", x"0080", x"0080", x"0080", x"0080", x"007F", x"007F", x"007F", x"007F", x"007E", x"007E", x"007E", x"007E", x"007D", x"007D", x"007D", x"007D", x"007C", x"007C", x"007C", x"007C", x"007B", x"007B", x"007B", x"007B", x"007A", x"007A", x"007A", x"007A", x"0079", x"0079", x"0079", x"0079", x"0078", x"0078", x"0078", x"0078", x"0077", x"0077", x"0077", x"0077", x"0076", x"0076", x"0076", x"0076", x"0075", x"0075", x"0075", x"0075", x"0074", x"0074", x"0074", x"0074", x"0073", x"0073", x"0073", x"0073", x"0072", x"0072", x"0072", x"0072", x"0071", x"0071", x"0071", x"0071", x"0070", x"0070", x"0070", x"0070", x"006F", x"006F", x"006F", x"006F", x"006E", x"006E", x"006E", x"006E", x"006D", x"006D", x"006D", x"006D", x"006C", x"006C", x"006C", x"006C", x"006B", x"006B", x"006B", x"006B", x"006A", x"006A", x"006A", x"006A", x"0069", x"0069", x"0069", x"0069", x"0069", x"0068", x"0068", x"0068", x"0068", x"0067", x"0067", x"0067", x"0067", x"0066", x"0066", x"0066", x"0066", x"0065", x"0065", x"0065", x"0065", x"0064", x"0064", x"0064", x"0064", x"0063", x"0063", x"0063", x"0063", x"0063", x"0062", x"0062", x"0062", x"0062", x"0061", x"0061", x"0061", x"0061", x"0060", x"0060", x"0060", x"0060", x"005F", x"005F", x"005F", x"005F", x"005F", x"005E", x"005E", x"005E", x"005E", x"005D", x"005D", x"005D", x"005D", x"005C", x"005C", x"005C", x"005C", x"005B", x"005B", x"005B", x"005B", x"005B", x"005A", x"005A", x"005A", x"005A", x"0059", x"0059", x"0059", x"0059", x"0059", x"0058", x"0058", x"0058", x"0058", x"0057", x"0057", x"0057", x"0057", x"0056", x"0056", x"0056", x"0056", x"0056", x"0055", x"0055", x"0055", x"0055", x"0054", x"0054", x"0054", x"0054", x"0054", x"0053", x"0053", x"0053", x"0053", x"0053", x"0052", x"0052", x"0052", x"0052", x"0051", x"0051", x"0051", x"0051", x"0051", x"0050", x"0050", x"0050", x"0050", x"004F", x"004F", x"004F", x"004F", x"004F", x"004E", x"004E", x"004E", x"004E", x"004E", x"004D", x"004D", x"004D", x"004D", x"004C", x"004C", x"004C", x"004C", x"004C", x"004B", x"004B", x"004B", x"004B", x"004B", x"004A", x"004A", x"004A", x"004A", x"004A", x"0049", x"0049", x"0049", x"0049", x"0049", x"0048", x"0048", x"0048", x"0048", x"0048", x"0047", x"0047", x"0047", x"0047", x"0047", x"0046", x"0046", x"0046", x"0046", x"0046", x"0045", x"0045", x"0045", x"0045", x"0045", x"0044", x"0044", x"0044", x"0044", x"0044", x"0043", x"0043", x"0043", x"0043", x"0043", x"0042", x"0042", x"0042", x"0042", x"0042", x"0041", x"0041", x"0041", x"0041", x"0041", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"003F", x"003F", x"003F", x"003F", x"003F", x"003E", x"003E", x"003E", x"003E", x"003E", x"003E", x"003D", x"003D", x"003D", x"003D", x"003D", x"003C", x"003C", x"003C", x"003C", x"003C", x"003C", x"003B", x"003B", x"003B", x"003B", x"003B", x"003A", x"003A", x"003A", x"003A", x"003A", x"003A", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0038", x"0038", x"0038", x"0038", x"0038", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"002F", x"002F", x"002F", x"002F", x"002F", x"002F", x"002E", x"002E", x"002E", x"002E", x"002E", x"002E", x"002E", x"002D", x"002D", x"002D", x"002D", x"002D", x"002D", x"002D", x"002C", x"002C", x"002C", x"002C", x"002C", x"002C", x"002C", x"002B", x"002B", x"002B", x"002B", x"002B", x"002B", x"002B", x"002A", x"002A", x"002A", x"002A", x"002A", x"002A", x"002A", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"001F", x"001F", x"001F", x"001F", x"001F", x"001F", x"001F", x"001F", x"001F", x"001E", x"001E", x"001E", x"001E", x"001E", x"001E", x"001E", x"001E", x"001E", x"001D", x"001D", x"001D", x"001D", x"001D", x"001D", x"001D", x"001D", x"001D", x"001D", x"001C", x"001C", x"001C", x"001C", x"001C", x"001C", x"001C", x"001C", x"001C", x"001C", x"001B", x"001B", x"001B", x"001B", x"001B", x"001B", x"001B", x"001B", x"001B", x"001B", x"001B", x"001A", x"001A", x"001A", x"001A", x"001A", x"001A", x"001A", x"001A", x"001A", x"001A", x"001A", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000F", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000E", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000D", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000C", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000B", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"000A", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000");
begin
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (en = '1') then
                dout <= lut(to_integer(signed(din) + 4096));
            end if;
        end if;
    end process;
end Behavioral;
